module system_ctrl_tb ();
//parameters

//stubs

//output

//instance

//sim flow

endmodule